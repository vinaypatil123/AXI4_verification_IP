`include "uvm_macros.svh"

package axi;
  `include "axi_master_sequence_item.sv"
  `include "axi_master_sequence.sv"
  `include "axi_master_sequencer.sv"
  `include "axi_master_driver.sv"
  `include "axi_master_monitor.sv"
  `include "axi_master_configuration.sv"
endpackage : axi