import uvm_pkg::*;
`include "uvm_macros.svh"

`include "axi_interface.sv"
`include "axi_master_sequence_item.sv"
`include "axi_master_sequence.sv"
`include "axi_master_sequencer.sv"
`include "axi_master_driver.sv"
`include "axi_master_monitor.sv"
`include "axi_master_configuration.sv"
`include "axi_master_agent.sv"
`include "axi_environment.sv"
`include "axi_test.sv"
`include "axi_top.sv"